module EX(

);

endmodule

// PC加法器
module ysyx_22040088_pc_adder(
    input       [63:0] in,
    output      [63:0] out
);

assign out = in + 4;

endmodule